library verilog;
use verilog.vl_types.all;
entity bemicro_tb is
end bemicro_tb;
